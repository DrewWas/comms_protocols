
module rx #(
    parameters
) (
    input logic clk,
    input logic reset,
    
);
    
endmodule




